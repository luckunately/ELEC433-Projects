module HammingIn (
    input logic [63:0] data_in,
    output logic [71:0] data_out,
    output logic resend
)


endmodule